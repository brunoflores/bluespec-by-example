function Word alu (Word a, Word b, AluFunc f);
function Bool aluBr (Word a, Word b, BrFunc f);
